.include osu018.lib
.include sub_ckts.lib

XX1 N001 N005 N002 VDD 0 nand201
XX2 N002 N008 N006 VDD 0 nand201
XX3 N006 N007 N008 VDD 0 nand201
XX4 N007 N010 N011 VDD 0 nand201
XX5 N011 N009 N010 VDD 0 nand201
XX6 N013 N012 N009 VDD 0 nand201
XX7 f_clk_in N005 VDD 0 inv101
XX8 f_VCO N013 VDD 0 inv101
XX9 N002 N003 VDD 0 inv101
XX10 N003 N004 VDD 0 inv101
XX11 N009 N014 VDD 0 inv101
XX12 N014 N015 VDD 0 inv101
XX13 N004 N006 N007 N001 VDD 0 nand301
XX14 N007 N010 N015 N012 VDD 0 nand301
XX15 N012 down VDD 0 inv101
XX16 N006 N002 N009 N010 N007 VDD 0 nand401
XX17 N001 up VDD 0 inv101

V1 f_clk_in 0 pulse 0 1.8 0 100p 100p 5n 10n
V2 f_VCO 0 pulse 0 1.8 2n 100p 100p 5n 9n
V3 VDD 0 1.8


.control
tran .1ns 50n
plot V(f_clk_in)+6 V(f_VCO)+4 V(up)+2 V(down)
.endc


.end
