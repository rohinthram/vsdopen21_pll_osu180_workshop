* PFD with charge pump
.include osu018.lib
.include sub_ckts.lib

XX1 f_in f_out_8 up down pfd_501
XX2 up down vin_vco charge_pump


*___________LPF________________*
C1 Vin_vco 0 200p
C2 N001 0 500p
R1 Vin_vco N001 500
*______________________________*

V1 f_in 0 PULSE 0 1.8 10p 60p 60p 100n 200n
V2 f_out_8 0 PULSE 0 1.8 40n 60p 60p 100n 180n
V3 VDD 0 1.8


.control
tran .1n 4u
plot V(f_in)+8 V(f_out_8)+6 V(up)+4 V(down)+2 V(vin_vco)
.endc


.end



.subckt pfd_501 f_clk_in f_VCO up down
XX1 N001 N005 N002 vddd 0 nand201
XX2 N002 N008 N006 vddd 0 nand201
XX3 N006 N007 N008 vddd 0 nand201
XX4 N007 N010 N011 vddd 0 nand201
XX5 N011 N009 N010 vddd 0 nand201
XX6 N013 N012 N009 vddd 0 nand201
XX7 f_clk_in N005 vddd 0 inv101
XX8 f_VCO N013 vddd 0 inv101
XX9 N002 N003 vddd 0 inv101
XX10 N003 N004 vddd 0 inv101
XX11 N009 N014 vddd 0 inv101
XX12 N014 N015 vddd 0 inv101
XX13 N004 N006 N007 N001 vddd 0 nand301
XX14 N007 N010 N015 N012 vddd 0 nand301
XX15 N012 down vddd 0 inv101
XX16 N006 N002 N009 N010 N007 vddd 0 nand401
XX17 N001 up vddd 0 inv101
V1 vddd 0 1.8
.ends pfd_501

.subckt charge_pump UP Down CP
M7 UP_bar UP 0 0 nfet l=180n w=180n
M8 DOWN_bar Down 0 0 nfet l=180n w=180n
M12 VDD Down DOWN_bar VDD pfet l=180n w=540n
M14 VDD UP UP_bar VDD pfet l=180n w=540n
M15 UP_bar 0 N001 N001 nfet l=180n w=180n
M16 DOWN_bar 0 N004 N004 nfet l=180n w=180n
M17 N003 N004 N003 N003 nfet l=180n w=180n
M18 0 VDD VDD 0 nfet l=180n w=180n
M19 CP VDD N003 N003 nfet l=180n w=180n
M20 N003 Down 0 0 nfet l=180n w=15u
M21 N001 VDD UP_bar N001 pfet l=180n w=540n
M22 N004 VDD DOWN_bar N004 pfet l=180n w=540n
M23 N002 UP N002 N002 pfet l=180n w=540n
M24 0 0 VDD VDD pfet l=180n w=540n
M25 N002 0 CP N002 pfet l=180n w=540n
M26 VDD N001 N002 VDD pfet l=180n w=45u
V4 VDD 0 1.8
.ends charge_pump
