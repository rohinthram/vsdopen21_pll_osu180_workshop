.include osu018.lib

M3  out201 in1 Net-_M3-Pad3_ gnd nfet l=180n w=720n		
M4  Net-_M3-Pad3_ in2 gnd gnd nfet l=180n w=720n
M2  vdd in2 out201 vdd pfet l=180n w=360n
M1  vdd in1 out201 vdd pfet l=180n w=360n


v1 vdd gnd 1.8
v2 in1 gnd PULSE(0 1.8 0 .1u .1u 1u 2u) 
v3 in2 gnd PULSE(0 1.8 .5u .1u .1u 1u 1.9u)


.tran 1us 10u
.control
run
plot v(in1)+4 V(in2)+2 v(out201)
.endc	

.end
