.include osu018.lib

M1  out in gnd gnd nfet l=180n w=180n		
M2  vdd in out vdd pfet l=180n w=360n

v1 vdd gnd 1.8
v2 in gnd PULSE(0 1.8 0 .1u .1u 1u 2u) 


.tran 1us 10u
.control
run
plot v(in)+3 v(out)
.endc		

.end
