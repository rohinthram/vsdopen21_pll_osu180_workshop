.include osu018.lib

M4  out301 in1 Net-_M4-Pad3_ gnd nfet l=180n w=720n		
M5  Net-_M4-Pad3_ in2 Net-_M5-Pad3_ gnd nfet l=180n w=720n		
M6  Net-_M5-Pad3_ in3 gnd gnd nfet l=180n w=720n		
M2  vdd in2 out301 vdd pfet l=180n w=360n		
M3  vdd in3 out301 vdd pfet l=180n w=360n		
M1  vdd in1 out301 vdd pfet l=180n w=360n

v1 vdd gnd 1.8
v2 in1 gnd PULSE(0 1.8 0 .1u .1u 1u 2u) 
v3 in2 gnd PULSE(0 1.8 .5u .1u .1u 1u 1.9u)
v4 in3 gnd PULSE(0 1.8 .5u .1u .1u 1u 2.1u)

.tran 1us 10u
.control
run
plot v(in1)+6 v(in2)+4 V(in3)+2 v(out301)
.endc		

.end
