* /home/rohinth/Desktop/esim_simulation/nand401/nand401.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: Tue Oct 19 15:42:42 2021

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
M1  vdd in1 out401 vdd mosfet_p		
M2  vdd in2 out401 vdd mosfet_p		
M7  vdd in3 out401 vdd mosfet_p		
M8  vdd in4 out401 vdd mosfet_p		
M3  out401 in1 Net-_M3-Pad3_ gnd mosfet_n		
M4  Net-_M3-Pad3_ in2 Net-_M4-Pad3_ gnd mosfet_n		
M5  Net-_M4-Pad3_ in3 Net-_M5-Pad3_ gnd mosfet_n		
M6  Net-_M5-Pad3_ in4 gnd gnd mosfet_n		

.end
